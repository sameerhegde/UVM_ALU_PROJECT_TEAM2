//------------------------------------------------------------------------------
// Project      : ALU 
// File Name    : alu_package.sv
// Developers   : Vinod (5289) 
// Created Date : 03/09/2024
// Version      : V1.0
//------------------------------------------------------------------------------
// Copyright    : 2024(c) Manipal Center of Excellence. All rights reserved.
//------------------------------------------------------------------------------

`include "alu_sequence_item.v"
`include "alu_sequence.sv"
`include "alu_sequencer.sv"
`include "alu_driver.sv"
`include "alu_monitor_write.sv"
`include "alu_monitor_read.sv"
`include "alu_agent_active.sv"
`include "alu_agent_passive.sv"
`include "alu_scoreboard.sv"
`include "alu_coverage.sv"
`include "alu_environment.sv"
`include "alu_test.sv"
