//------------------------------------------------------------------------------
// Project      : ALU 
// File Name    : alu_define.svh
// Developers   : Team-2
// Created Date : 01/08/2024
// Version      : V1.0
//------------------------------------------------------------------------------
// Copyright    : 2024(c) Manipal Center of Excellence. All rights reserved.
//------------------------------------------------------------------------------

`timescale 10ns/100ps //Time Unit (ns) / Precision(ps)
`define WIDTH 8
`define NUM_TRANSACTIONS 4
`define CMD_WIDTH 4
