class alu_seq extends uvm_sequence #(alu_seq_item);

  // Factory registration
  `uvm_object_utils (alu_seq)

  // Class constructor
  function new (string name = "alu_seq");
    super.new (name);
  endfunction: new

  // Handle for alu_seq_item
  alu_seq_item txn;

  virtual task body;
    //repeat (`NUM_TRANSACTIONS) begin
      `uvm_info("SEQUENCE","start",UVM_LOW)
      txn = alu_seq_item::type_id::create("txn");
      wait_for_grant ();
      txn.randomize();
      send_request (txn);
      wait_for_item_done ();
    //end
  endtask: body

endclass: alu_seq

//-----------------------------------------------------------------------------
// ARITHMETIC OPERATIONS
//-----------------------------------------------------------------------------

// class alu_add_sequence extends uvm_sequence #(alu_seq_item);

//   `uvm_object_utils(alu_add_sequence)

//   function new(string name = "alu_add_sequence");
//     super.new(name);
//   endfunction
  
//   alu_seq_item txn;

//   virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//     txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0000; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//     if(txn.inp_valid == 2'b01 || txn.inp_valid == 2'b10) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//        txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0000;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//       txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0000;txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//   endtask
 
// endclass
//-------------------------------------------------------------------------------

class alu_sub_sequence extends uvm_sequence #(alu_seq_item);

  `uvm_object_utils(alu_sub_sequence)

  function new(string name = "alu_sub_sequence");
    super.new(name);
  endfunction
  
  alu_seq_item txn;

  virtual task body();
    txn = alu_seq_item::type_id::create("txn");
    wait_for_grant();
    txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0001; txn.delay < 8;txn.opa>txn.opb;};
    send_request(txn);
    wait_for_item_done();
   
    if(txn.inp_valid == 2'b01 || txn.inp_valid == 2'b10) begin
     txn.opa.rand_mode(0); 
     txn.opb.rand_mode(0);
     txn.inp_valid.rand_mode(0);
     txn.delay.rand_mode(0);
      repeat (txn.delay) begin
       txn.delay.rand_mode(0);
       wait_for_grant();
        txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0001;};
       send_request(txn);
       wait_for_item_done();
       end
      txn.inp_valid.rand_mode(1);
      //txn.delay.rand_mode(1);
      wait_for_grant();
      txn.randomize() with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0001;txn.inp_valid==2'b11;};
       send_request(txn);
       wait_for_item_done();
    end
  endtask
endclass
// //-------------------------------------------------------------------------------------
// class alu_add_cin_seq extends alu_seq;

//   `uvm_object_utils(alu_add_cin_seq)

//   function new(string name = "alu_add_cin_seq");
//     super.new(name);
//   endfunction

   
//   alu_seq_item txn;

//   virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//     txn.randomize()with {txn.mode == 1; txn.ce == 1;txn.cin == 1; txn.cmd == 4'b0010; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//     if(txn.inp_valid == 2'b01 || txn.inp_valid == 2'b10) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//         txn.randomize()with {txn.mode == 1; txn.ce == 1;txn.cin == 1; txn.cmd == 4'b0010;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//       txn.randomize()with {txn.mode == 1; txn.ce == 1;txn.cin == 1; txn.cmd == 4'b0010;txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//   endtask
// endclass
//-------------------------------------------------------------------------------------------------------
// class alu_sub_cin_seq extends alu_seq;

//   `uvm_object_utils(alu_sub_cin_seq)

//   function new(string name = "alu_sub_cin_seq");
//     super.new(name);
//   endfunction
 
//   alu_seq_item txn;

//   virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//     txn.randomize()with {txn.mode == 1; txn.ce == 1;txn.cin == 1; txn.cmd == 4'b0011; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//     if(txn.inp_valid == 2'b01 || txn.inp_valid == 2'b10) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//         txn.randomize()with {txn.mode == 1; txn.ce == 1;txn.cin == 1; txn.cmd == 4'b0011;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//       txn.randomize()with {txn.mode == 1; txn.ce == 1;txn.cin == 1; txn.cmd == 4'b0011;txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//   endtask
// endclass

//---------------------------------------------------------------------------------------------------

class alu_inc_opa_seq extends alu_seq;

  `uvm_object_utils(alu_inc_opa_seq)

  function new(string name = "alu_inc_opa_seq");
    super.new(name);
  endfunction

 alu_seq_item txn;

  virtual task body();
    txn = alu_seq_item::type_id::create("txn");
    wait_for_grant();
    txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0100; txn.delay < 8;};
    send_request(txn);
    wait_for_item_done();
   
    if(txn.inp_valid == 2'b10) begin
     txn.opa.rand_mode(0); 
     txn.opb.rand_mode(0);
     txn.inp_valid.rand_mode(0);
     txn.delay.rand_mode(0);
      repeat (txn.delay) begin
       txn.delay.rand_mode(0);
       wait_for_grant();
        txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0100;};
       send_request(txn);
       wait_for_item_done();
       end
      txn.inp_valid.rand_mode(1);
      //txn.delay.rand_mode(1);
      wait_for_grant();
      txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0100;txn.inp_valid==2'b01||txn.inp_valid==2'b11;};
       send_request(txn);
       wait_for_item_done();
    end
    endtask
endclass

// //-------------------------------------------------------------------------------------------
// class alu_dec_opa_seq extends alu_seq;

//   `uvm_object_utils(alu_dec_opa_seq)

//   function new(string name = "alu_dec_opa_seq");
//     super.new(name);
//   endfunction
//   alu_seq_item txn;

//  virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//    txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0101; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//     if(txn.inp_valid == 2'b10) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//         txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0101;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//       txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0101;txn.inp_valid==2'b01;txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//     endtask
// endclass
// //--------------------------------------------------------------------------------------------------------
// class alu_inc_opb_seq extends alu_seq;

//   `uvm_object_utils(alu_inc_opb_seq)

//   function new(string name = "alu_inc_opb_seq");
//     super.new(name);
//   endfunction
// alu_seq_item txn;

//  virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//    txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0110; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//    if(txn.inp_valid == 2'b01) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//         txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0110;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//       txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0110;txn.inp_valid==2'b10;txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//     endtask
// endclass

// //-------------------------------------------------------------------------------------------------
// class alu_dec_opb_seq extends alu_seq;

//   `uvm_object_utils(alu_dec_opb_seq)

//   function new(string name = "alu_dec_opb_seq");
//     super.new(name);
//   endfunction
// alu_seq_item txn;

//  virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//    txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0111; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//    if(txn.inp_valid == 2'b01) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//         txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0111;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//      txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b0111;txn.inp_valid==2'b10;txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//     endtask
// endclass
// //-----------------------------------------------------------------------------------------
// class alu_cmp_seq extends alu_seq;

//   `uvm_object_utils(alu_cmp_seq)

//   function new(string name = "alu_cmp_seq");
//     super.new(name);
//   endfunction
//   alu_seq_item txn;
//  virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//    txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1000; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//    if(txn.inp_valid == 2'b01 || txn.inp_valid ==2'b10) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//         txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1000;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//      txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1000; txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//     endtask
// endclass

// //---------------------------------------------------------------------------------------------------
// class alu_inc_mul_seq extends alu_seq;

//   `uvm_object_utils(alu_inc_mul_seq)

//   function new(string name = "alu_inc_mul_seq");
//     super.new(name);
//   endfunction
  
//  alu_seq_item txn;
  
//  virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//    txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1001; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//    if(txn.inp_valid == 2'b01 || txn.inp_valid ==2'b10) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//         txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1001;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//      txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1001; txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//     endtask
// endclass
// //---------------------------------------------------------------------------------------------
// class alu_opa_lshift_mul_seq extends alu_seq;

//   `uvm_object_utils(alu_opa_lshift_mul_seq)

//   function new(string name = "alu_opa_lshift_mul_seq");
//     super.new(name);
//   endfunction
  
//  alu_seq_item txn;
  
//   virtual task body();
//     txn = alu_seq_item::type_id::create("txn");
//     wait_for_grant();
//     txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1010; txn.delay < 8;};
//     send_request(txn);
//     wait_for_item_done();
   
//    if(txn.inp_valid == 2'b01 || txn.inp_valid ==2'b10) begin
//      txn.opa.rand_mode(0); 
//      txn.opb.rand_mode(0);
//      txn.inp_valid.rand_mode(0);
//      txn.delay.rand_mode(0);
//       repeat (txn.delay) begin
//        txn.delay.rand_mode(0);
//        wait_for_grant();
//         txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1010;};
//        send_request(txn);
//        wait_for_item_done();
//        end
//       txn.inp_valid.rand_mode(1);
//       //txn.delay.rand_mode(1);
//       wait_for_grant();
//      txn.randomize()with {txn.mode == 1; txn.ce == 1; txn.cmd == 4'b1010; txn.inp_valid==2'b11;};
//        send_request(txn);
//        wait_for_item_done();
//     end
//     endtask
// endclass
// //----------------------------------------------------------------------------------x	


